library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package platform_variant_pkg is


-- Super Earth Invasion
	constant ROM_0_NAME		: string := "roms/searthin.hex";
	constant ROM_1_NAME		: string := "";
	constant VRAM_NAME		: string := "";
end;